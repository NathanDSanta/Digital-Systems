LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY MUX4 IS
  PORT (
    SEL        : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    A, B, C, D : IN STD_LOGIC;
    F          : OUT STD_LOGIC);
END MUX;
ARCHITECTURE BEHAVIOUR OF MUX4 IS
  SIGNAL SEL1, SEL1B, SEL0, SEL0B;
BEGIN
  SEL1  <= SEL(1);
  SEL1B <= NOT SEL(1);
  SEL0  <= SEL(0);
  SEL0B <= NOT SEL(0);
  F     <= (A AND SEL1B AND SEL0B) OR
  (B AND SEL1B AND SEL0) OR
  (C AND SEL1 AND SEL0B) OR
  (D AND SEL1 AND SEL0);
END;
